magic
tech sky130A
magscale 1 2
timestamp 1729223408
<< nwell >>
rect -203 -633 997 565
<< nsubdiff >>
rect -167 495 -107 529
rect 901 495 961 529
rect -167 469 -133 495
rect 927 469 961 495
rect -167 -563 -133 -537
rect 927 -563 961 -537
rect -167 -597 -107 -563
rect 901 -597 961 -563
<< nsubdiffcont >>
rect -107 495 901 529
rect -167 -537 -133 469
rect 927 -537 961 469
rect -107 -597 901 -563
<< poly >>
rect -40 397 48 413
rect -40 363 -24 397
rect 10 363 48 397
rect -40 342 48 363
rect 738 397 814 413
rect 738 363 764 397
rect 798 363 814 397
rect 738 341 814 363
rect -43 -428 48 -404
rect -43 -462 -27 -428
rect 7 -462 48 -428
rect -43 -478 48 -462
rect 738 -428 826 -407
rect 738 -462 776 -428
rect 810 -462 826 -428
rect 738 -478 826 -462
<< polycont >>
rect -24 363 10 397
rect 764 363 798 397
rect -27 -462 7 -428
rect 776 -462 810 -428
<< locali >>
rect -167 495 -107 529
rect 901 495 961 529
rect -167 469 -133 495
rect 927 469 961 495
rect -40 363 -24 397
rect 10 363 26 397
rect 748 363 764 397
rect 798 363 814 397
rect -43 -462 -27 -428
rect 7 -462 23 -428
rect 760 -462 776 -428
rect 810 -462 826 -428
rect -167 -563 -133 -537
rect 927 -563 961 -537
rect -167 -597 -107 -563
rect 901 -597 961 -563
<< viali >>
rect -24 363 10 397
rect 764 363 798 397
rect -27 -462 7 -428
rect 776 -462 810 -428
<< metal1 >>
rect -100 431 892 464
rect -100 -496 -67 431
rect -36 397 22 403
rect -36 363 -24 397
rect 10 363 22 397
rect -36 357 22 363
rect -27 307 6 357
rect 124 333 188 403
rect 282 397 346 403
rect 376 397 409 431
rect 440 397 504 403
rect 282 364 504 397
rect 282 333 346 364
rect 440 333 504 364
rect 598 333 662 403
rect 752 397 810 403
rect 752 363 764 397
rect 798 363 820 397
rect 752 357 820 363
rect 780 304 820 357
rect -28 180 94 304
rect 692 292 820 304
rect 692 180 814 292
rect -28 128 42 180
rect 94 128 104 180
rect 199 128 209 180
rect 261 128 271 180
rect -39 69 15 79
rect 124 69 188 98
rect 13 35 188 69
rect 13 17 22 35
rect 124 28 188 35
rect 282 29 346 99
rect -39 7 15 17
rect 376 -4 410 131
rect 515 128 525 180
rect 577 128 587 180
rect 682 128 692 180
rect 744 128 814 180
rect 440 28 504 98
rect 598 69 662 99
rect 764 69 826 79
rect 598 35 774 69
rect 598 29 662 35
rect 764 17 774 35
rect 764 7 826 17
rect 57 -38 726 -4
rect 57 -193 91 -38
rect 124 -164 188 -94
rect 282 -100 346 -94
rect 440 -100 504 -94
rect 278 -152 288 -100
rect 340 -134 446 -100
rect 340 -152 350 -134
rect 436 -152 446 -134
rect 498 -152 508 -100
rect 282 -164 346 -152
rect 440 -164 504 -152
rect 598 -164 662 -94
rect 692 -193 726 -38
rect -31 -369 91 -193
rect 199 -245 209 -193
rect 261 -245 271 -193
rect 357 -245 367 -193
rect 419 -245 429 -193
rect 515 -245 525 -193
rect 577 -245 587 -193
rect 689 -220 811 -193
rect 690 -225 811 -220
rect 689 -364 811 -225
rect 689 -369 814 -364
rect -28 -422 7 -369
rect -39 -428 19 -422
rect -39 -462 -27 -428
rect 7 -462 19 -428
rect -39 -468 19 -462
rect 124 -468 188 -398
rect 282 -468 346 -398
rect 440 -468 504 -398
rect 598 -468 662 -398
rect 780 -422 814 -369
rect 764 -428 822 -422
rect 764 -462 776 -428
rect 810 -462 822 -428
rect 764 -468 822 -462
rect 139 -496 172 -468
rect 613 -496 646 -468
rect 859 -496 892 431
rect -100 -529 892 -496
<< via1 >>
rect 42 128 94 180
rect 209 128 261 180
rect -39 17 13 69
rect 525 128 577 180
rect 692 128 744 180
rect 774 17 826 69
rect 288 -152 340 -100
rect 446 -152 498 -100
rect 209 -245 261 -193
rect 367 -245 419 -193
rect 525 -245 577 -193
<< metal2 >>
rect 218 194 252 207
rect 42 180 94 190
rect 42 116 94 128
rect 207 184 263 194
rect 207 118 263 128
rect 523 184 579 194
rect 523 118 579 128
rect 692 180 744 190
rect 692 118 744 128
rect -40 69 13 79
rect -40 17 -39 69
rect -40 7 13 17
rect -30 -100 2 7
rect 42 -2 86 116
rect 700 -2 744 118
rect 774 69 826 79
rect 774 7 826 17
rect 42 -46 744 -2
rect 288 -100 340 -90
rect -30 -134 288 -100
rect 288 -162 340 -152
rect 371 -183 415 -46
rect 446 -100 498 -90
rect 784 -100 816 7
rect 498 -134 816 -100
rect 446 -162 498 -152
rect 207 -193 263 -183
rect 207 -259 263 -249
rect 367 -193 419 -183
rect 367 -255 419 -245
rect 523 -193 579 -183
rect 523 -259 579 -249
<< via2 >>
rect 207 180 263 184
rect 207 128 209 180
rect 209 128 261 180
rect 261 128 263 180
rect 523 180 579 184
rect 523 128 525 180
rect 525 128 577 180
rect 577 128 579 180
rect 207 -245 209 -193
rect 209 -245 261 -193
rect 261 -245 263 -193
rect 207 -249 263 -245
rect 523 -245 525 -193
rect 525 -245 577 -193
rect 577 -245 579 -193
rect 523 -249 579 -245
<< metal3 >>
rect 197 184 273 253
rect 197 128 207 184
rect 263 128 273 184
rect 197 123 273 128
rect 513 184 589 253
rect 513 128 523 184
rect 579 128 589 184
rect 513 123 589 128
rect 204 -26 266 123
rect 523 -26 585 123
rect 204 -88 585 -26
rect 204 -188 266 -88
rect 523 -188 585 -88
rect 197 -193 273 -188
rect 197 -249 207 -193
rect 263 -249 273 -193
rect 197 -318 273 -249
rect 513 -193 589 -188
rect 513 -249 523 -193
rect 579 -249 589 -193
rect 513 -318 589 -249
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729183152
transform 1 0 753 0 1 -281
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729183152
transform 1 0 753 0 1 216
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729183152
transform 1 0 33 0 1 216
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729183152
transform 1 0 33 0 1 -281
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_V8EW6L  sky130_fd_pr__pfet_01v8_V8EW6L_0
timestamp 1729183152
transform 1 0 393 0 1 216
box -381 -200 381 200
use sky130_fd_pr__pfet_01v8_V8EW6L  sky130_fd_pr__pfet_01v8_V8EW6L_1
timestamp 1729183152
transform 1 0 393 0 1 -281
box -381 -200 381 200
<< labels >>
flabel nsubdiffcont 391 507 391 507 0 FreeSans 480 0 0 0 VDD
port 0 nsew
flabel via1 75 151 75 151 0 FreeSans 480 0 0 0 D6
port 1 nsew
flabel via2 232 147 232 147 0 FreeSans 480 0 0 0 S67
port 2 nsew
flabel via1 -16 46 -16 46 0 FreeSans 480 0 0 0 VIN
port 3 nsew
flabel metal1 61 -272 61 -272 0 FreeSans 480 0 0 0 OUT
port 4 nsew
flabel metal1 159 -451 159 -451 0 FreeSans 480 0 0 0 VIP
port 5 nsew
<< end >>

** sch_path: /home/surya/Ring_Oscilator/ring_oscillator.sch
**.subckt ring_oscillator vdd out gnd
*.iopin vdd
*.iopin gnd
*.opin out
x1 vdd out net1 gnd inverter
x2 vdd net1 net2 gnd inverter
x3 vdd net2 out gnd inverter
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/surya/Ring_Oscilator/inverter.sym
** sch_path: /home/surya/Ring_Oscilator/inverter.sch

.end

magic
tech sky130A
magscale 1 2
timestamp 1729053250
<< metal1 >>
rect 296 2380 1670 2512
rect 398 2108 442 2380
rect 822 2104 866 2380
rect 1244 2104 1288 2380
rect 502 1914 564 1920
rect 502 1858 508 1914
rect 560 1858 564 1914
rect 1494 1914 1632 1920
rect 652 1872 1020 1904
rect 1072 1870 1440 1902
rect 502 1850 564 1858
rect 1494 1862 1510 1914
rect 1614 1862 1632 1914
rect 1494 1850 1632 1862
rect 402 1398 446 1668
rect 824 1398 868 1668
rect 1246 1398 1290 1672
rect 298 1266 1672 1398
<< via1 >>
rect 508 1858 560 1914
rect 1510 1862 1614 1914
<< metal2 >>
rect 502 1914 1632 1920
rect 502 1858 508 1914
rect 560 1862 1510 1914
rect 1614 1862 1632 1914
rect 560 1858 1632 1862
rect 502 1850 1632 1858
use inverter  x1
timestamp 1728978940
transform 1 0 423 0 1 1306
box -53 21 369 1147
use inverter  x2
timestamp 1728978940
transform 1 0 844 0 1 1306
box -53 21 369 1147
use inverter  x3
timestamp 1728978940
transform 1 0 1265 0 1 1306
box -53 21 369 1147
<< labels >>
flabel metal1 308 2486 308 2486 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel metal2 1626 1884 1626 1884 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 346 1302 346 1302 0 FreeSans 320 0 0 0 GND
port 3 nsew
<< end >>

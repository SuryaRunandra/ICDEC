magic
tech sky130A
magscale 1 2
timestamp 1728974160
<< checkpaint >>
rect -1260 -1260 2051 2766
use untitled-1  x1
timestamp 1728974159
transform 1 0 53 0 1 1306
box -53 -1306 738 200
<< end >>

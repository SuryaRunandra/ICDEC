magic
tech sky130A
magscale 1 2
timestamp 1729415910
<< metal1 >>
rect 3190 2652 3220 2680
rect 241 1774 251 1826
rect 303 1774 313 1826
rect 1404 1768 1414 1820
rect 1466 1768 1476 1820
rect 1543 1613 1583 1647
rect 1640 1355 1674 1389
rect 2170 1367 2574 1401
rect 1865 1265 1875 1317
rect 1927 1265 1937 1317
rect 2170 1308 2204 1367
rect 2540 1253 2574 1367
rect 1755 968 1787 1017
<< via1 >>
rect 251 1774 303 1826
rect 1414 1768 1466 1820
rect 1875 1265 1927 1317
<< metal2 >>
rect 255 2211 1491 2254
rect 255 1836 298 2211
rect 1378 2105 1409 2144
rect 251 1826 303 1836
rect 1414 1820 1466 1830
rect 251 1764 303 1774
rect 786 1780 1414 1810
rect 786 1697 816 1780
rect 1414 1758 1466 1768
rect 1885 1436 2589 1468
rect 1885 1327 1917 1436
rect 1875 1317 1927 1327
rect 1875 1255 1927 1265
<< metal3 >>
rect 1930 2310 2616 2372
rect 1930 2239 1992 2310
use nmosamp  nmosamp_0
timestamp 1729221421
transform 1 0 292 0 1 1074
box -292 -1074 733 955
use nmoscs  nmoscs_0
timestamp 1729173886
transform 1 0 1370 0 1 748
box -346 -748 1034 694
use pmosamp  pmosamp_0
timestamp 1729223408
transform 1 0 1407 0 1 2075
box -203 -633 997 565
use pmoscs  pmoscs_0
timestamp 1729152682
transform 1 0 2584 0 1 1461
box -180 -1461 818 1419
<< labels >>
flabel metal2 1088 1792 1088 1792 0 FreeSans 2080 0 0 0 OUT
port 0 nsew
flabel metal1 3204 2658 3204 2658 0 FreeSans 2080 0 0 0 VDD
port 1 nsew
flabel metal1 1659 1372 1659 1372 0 FreeSans 2080 0 0 0 GND
port 2 nsew
flabel metal2 1389 2123 1389 2123 0 FreeSans 2080 0 0 0 VIN
port 3 nsew
flabel metal1 1563 1630 1563 1630 0 FreeSans 2080 0 0 0 VIP
port 4 nsew
flabel metal1 1773 991 1773 991 0 FreeSans 2080 0 0 0 RS
port 5 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1728974159
<< checkpaint >>
rect -944 -2566 1998 574
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 0
transform 1 0 158 0 1 -934
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 0
transform 1 0 527 0 1 -996
box -211 -310 211 310
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 out
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 gnd
port 3 nsew
<< end >>

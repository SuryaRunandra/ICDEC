magic
tech sky130A
magscale 1 2
timestamp 1728978907
<< viali >>
rect 57 202 91 378
rect 57 -428 91 -252
<< metal1 >>
rect 51 378 190 390
rect 51 202 57 378
rect 91 202 190 378
rect 51 190 190 202
rect 257 190 369 253
rect 215 -202 249 143
rect 306 -240 369 190
rect 51 -252 188 -240
rect 51 -428 57 -252
rect 91 -428 189 -252
rect 253 -303 369 -240
rect 51 -440 97 -428
use sky130_fd_pr__pfet_01v8_LGS3BL  XM1
timestamp 1728978907
transform 1 0 232 0 1 254
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM2
timestamp 1728978907
transform 1 0 232 0 1 -309
box -211 -279 211 279
<< labels >>
flabel metal1 133 267 133 267 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 127 -337 127 -337 0 FreeSans 160 0 0 0 GND
port 2 nsew
flabel metal1 338 -26 338 -26 0 FreeSans 160 0 0 0 OUT
port 3 nsew
flabel metal1 233 -31 233 -31 0 FreeSans 160 0 0 0 IN
port 4 nsew
<< end >>
